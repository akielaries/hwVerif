module top;
    initial begin
        $display("Hello World!");
        $finish;
    end
endmodule


