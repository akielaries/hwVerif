module two_bit_comp(
    input [1:0] input_a,
    input [1:0] input_b,
    output output_a
    );



endmodule

