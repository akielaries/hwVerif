/*
 * 2-bit comparator
 *
 * RANGE : 
 *      0 TO 2^n - 1
 *      0 TO 2^2 - 1 = 3
 *      0 TO 3
 */

module two_bit_comp(
    input [1:0] input_a,
    input [1:0] input_b,
    output output_a
    );



endmodule

