module hello;
    initial begin
        $display("Hello via verilog");
        $finish;
    end
endmodule

